module regfile (input  logic clk, we3,
                input  logic [4:0] ra1, ra2, wa3,
                input  logic [63:0] wd3,
                output logic [64:0] rd1, rd2);

    /*Banco de registros*/
endmodule